library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pong_game_over is 
    port(
        pixel_x : in STD_LOGIC_VECTOR (9 downto 0);
        pixel_y : in STD_LOGIC_VECTOR (9 downto 0);
        life_cnt: in STD_LOGIC_VECTOR (1 downto 0);
        game_over_on: out std_logic;
        graph_rgb: out std_logic_vector(2 downto 0)
    );
end pong_game_over;

architecture arch of pong_game_over is 
    -- x, y coordinates (0,0 to (639, 479)
    signal pix_x, pix_y: unsigned(9 downto 0);
    signal char_rgb: std_logic_vector (2 downto 0);
    -- screen dimensions
    constant MAX_X: integer := 640;
    constant MAX_Y: integer := 480;

    signal life_cnter: unsigned (1 downto 0);

    constant CHAR_SIZE: integer := 50;
    type char_type is array (0 to 49) of std_logic_vector (0 to 49);
    constant U_ROM: char_type := (
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "11111100000000000000000000000000000000000011111100",
        "01111110000000000000000000000000000000000111111000",
        "00111111000000000000000000000000000000001111110000",
        "00011111100000000000000000000000000000011111100000",
        "00001111110000000000000000000000000000111111000000",
        "00000111111111111111111111111111111111111110000000",
        "00000011111111111111111111111111111111111100000000",
        "00000001111111111111111111111111111111111000000000"
    );
    constant D_1_ROM: char_type := (
        "00000000000000000000000000000000000011111111111111",
        "00000000000000000000000000000000011111111111111111",
        "00000000000000000000000000000011111111111111111111",
        "00000000000000000000000000011111111111111111111111",
        "00000000000000000000000011111111111111111111111111",
        "00000000000000000000001111111111111111111111111111",
        "00000000000000000000111111111111111111111111111111",
        "00000000000000000011111111111111111111111111111111",
        "00000000000000001111111111111111111111111111111111",
        "00000000000000111111111111111111111111111111111111",
        "00000000000011111111111111111111111111111111111111",
        "00000000111111111111111111111111111111111111111111",
        "00000011111111111111111111111111111111111111111111",
        "00001111111111111111111111111111111111111111111111",
        "00011111111111111111111111111111111111111111111111",
        "00111111111111111111111111111111111111111111111111",
        "01111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111111111111111111111111111111111111",
        "01111111111111111111111111111111111111111111111111",
        "00111111111111111111111111111111111111111111111111",
        "00011111111111111111111111111111111111111111111111",
        "00001111111111111111111111111111111111111111111111",
        "00000111111111111111111111111111111111111111111111",
        "00000011111111111111111111111111111111111111111111",
        "00000001111111111111111111111111111111111111111111",
        "00000000111111111111111111111111111111111111111111",
        "00000000011111111111111111111111111111111111111111",
        "00000000001111111111111111111111111111111111111111",
        "00000000000111111111111111111111111111111111111111",
        "00000000000011111111111111111111111111111111111111",
        "00000000000000111111111111111111111111111111111111"
    );
    constant I_ROM: char_type := (
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "00000000000000000000111111111100000000000000000000",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111"
    );
    constant E_ROM: char_type := (
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "00000000000000000000000000000000000000000000011111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111"
    );
    constant D_2_ROM: char_type := (
        "00000000000000000000000000000000000011111111111111",
        "00000000000000000000000000000000011111111111111111",
        "00000000000000000000000000000011111111111111111111",
        "00000000000000000000000000011111111111111111111111",
        "00000000000000000000000011111111111111111111111111",
        "00000000000000000000001111111111111111111111111111",
        "00000000000000000000111111111111111111111111111111",
        "00000000000000000011111111111111111111111111111111",
        "00000000000000001111111111111111111111111111111111",
        "00000000000000111111111111111111111111111111111111",
        "00000000000011111111111111111111111111111111111111",
        "00000000111111111111111111111111111111111111111111",
        "00000011111111111111111111111111111111111111111111",
        "00001111111111111111111111111111111111111111111111",
        "00011111111111111111111111111111111111111111111111",
        "00111111111111111111111111111111111111111111111111",
        "01111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111111111111111111111111111111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111000000000000000000000011111111111",
        "11111111111111111111111111111111111111111111111111",
        "01111111111111111111111111111111111111111111111111",
        "00111111111111111111111111111111111111111111111111",
        "00011111111111111111111111111111111111111111111111",
        "00001111111111111111111111111111111111111111111111",
        "00000111111111111111111111111111111111111111111111",
        "00000011111111111111111111111111111111111111111111",
        "00000001111111111111111111111111111111111111111111",
        "00000000111111111111111111111111111111111111111111",
        "00000000011111111111111111111111111111111111111111",
        "00000000001111111111111111111111111111111111111111",
        "00000000000111111111111111111111111111111111111111",
        "00000000000011111111111111111111111111111111111111",
        "00000000000000111111111111111111111111111111111111"
    );

    constant U_X_L: integer := (MAX_X/2) - (CHAR_SIZE/2) - 1;
    constant U_X_R: integer:= U_X_L + CHAR_SIZE - 1;
    constant U_Y_T: integer := (MAX_Y/2) - (CHAR_SIZE/2) - 50;
    constant U_Y_B: integer:= U_Y_T + CHAR_SIZE - 1;

    constant D_1_X_L: integer := (MAX_X/2) - (4*(CHAR_SIZE/2)) - 1;
    constant D_1_X_R: integer:= D_1_X_L + CHAR_SIZE - 1;
    constant D_1_Y_T: integer := (MAX_Y/2) + (CHAR_SIZE/2) - 1;
    constant D_1_Y_B: integer:= D_1_Y_T + CHAR_SIZE - 1;

    constant I_X_L: integer := (MAX_X/2) - (2*(CHAR_SIZE/2)) - 1;
    constant I_X_R: integer:= I_X_L + CHAR_SIZE - 1;
    constant I_Y_T: integer := (MAX_Y/2) + (CHAR_SIZE/2) - 1;
    constant I_Y_B: integer:= I_Y_T + CHAR_SIZE - 1;

    constant E_X_L: integer := (MAX_X/2) + ((CHAR_SIZE/2)) - 1;
    constant E_X_R: integer:= E_X_L + CHAR_SIZE - 1;
    constant E_Y_T: integer := (MAX_Y/2) + (CHAR_SIZE/2) - 1;
    constant E_Y_B: integer:= E_Y_T + CHAR_SIZE - 1;

    constant D_2_X_L: integer := (MAX_X/2) + (4*(CHAR_SIZE/2)) - 1;
    constant D_2_X_R: integer:= D_2_X_L + CHAR_SIZE - 1;
    constant D_2_Y_T: integer := (MAX_Y/2) + (CHAR_SIZE/2) - 1;
    constant D_2_Y_B: integer:= D_2_Y_T + CHAR_SIZE - 1;

    signal rom_addr_U, rom_col_U: unsigned(5 downto 0);
    signal rom_data_U: std_logic_vector(49 downto 0);
    signal rom_bit_U: std_logic;
    signal sq_U_on: std_logic;
    signal U_cur_val_on: std_logic;
    signal U_y_t_u: unsigned(9 downto 0);
    signal U_x_l_u: unsigned(9 downto 0);

    signal rom_addr_D_1, rom_col_D_1: unsigned(5 downto 0);
    signal rom_data_D_1: std_logic_vector(49 downto 0);
    signal rom_bit_D_1: std_logic;
    signal sq_D_1_on: std_logic;
    signal D_1_cur_val_on: std_logic;
    signal D_1_y_t_u: unsigned(9 downto 0);
    signal D_1_x_l_u: unsigned(9 downto 0);

    signal rom_addr_I, rom_col_I: unsigned(5 downto 0);
    signal rom_data_I: std_logic_vector(49 downto 0);
    signal rom_bit_I: std_logic;
    signal sq_I_on: std_logic;
    signal I_cur_val_on: std_logic;
    signal I_y_t_u: unsigned(9 downto 0);
    signal I_x_l_u: unsigned(9 downto 0);

    signal rom_addr_E, rom_col_E: unsigned(5 downto 0);
    signal rom_data_E: std_logic_vector(49 downto 0);
    signal rom_bit_E: std_logic;
    signal sq_E_on: std_logic;
    signal E_cur_val_on: std_logic;
    signal E_y_t_u: unsigned(9 downto 0);
    signal E_x_l_u: unsigned(9 downto 0);

    signal rom_addr_D_2, rom_col_D_2: unsigned(5 downto 0);
    signal rom_data_D_2: std_logic_vector(49 downto 0);
    signal rom_bit_D_2: std_logic;
    signal sq_D_2_on: std_logic;
    signal D_2_cur_val_on: std_logic;
    signal D_2_y_t_u: unsigned(9 downto 0);
    signal D_2_x_l_u: unsigned(9 downto 0);

begin
    char_rgb <= "110"; -- red color characters

    pix_x <= unsigned(pixel_x);
    pix_y <= unsigned(pixel_y);
    life_cnter <= unsigned(life_cnt);

    sq_U_on <= '1' when (U_X_L <= pix_x) and (pix_x <= U_X_R) and (U_Y_T <= pix_y) and (pix_y <= U_Y_B) else '0';
    sq_D_1_on <= '1' when (D_1_X_L <= pix_x) and (pix_x <= D_1_X_R) and (D_1_Y_T <= pix_y) and (pix_y <= D_1_Y_B) else '0';
    sq_I_on <= '1' when (I_X_L <= pix_x) and (pix_x <= I_X_R) and (I_Y_T <= pix_y) and (pix_y <= I_Y_B) else '0';
    sq_E_on <= '1' when (E_X_L <= pix_x) and (pix_x <= E_X_R) and (E_Y_T <= pix_y) and (pix_y <= E_Y_B) else '0';
    sq_D_2_on <= '1' when (D_2_X_L <= pix_x) and (pix_x <= D_2_X_R) and (D_2_Y_T <= pix_y) and (pix_y <= D_2_Y_B) else '0';

    U_y_t_u <= to_unsigned(U_Y_T, 10);
    U_x_l_u <= to_unsigned(U_X_L, 10);

    D_1_y_t_u <= to_unsigned(D_1_Y_T, 10);
    D_1_x_l_u <= to_unsigned(D_1_X_L, 10);

    I_y_t_u <= to_unsigned(I_Y_T, 10);
    I_x_l_u <= to_unsigned(I_X_L, 10);

    E_y_t_u <= to_unsigned(E_Y_T, 10);
    E_x_l_u <= to_unsigned(E_X_L, 10);

    D_2_y_t_u <= to_unsigned(D_2_Y_T, 10);
    D_2_x_l_u <= to_unsigned(D_2_X_L, 10);

    rom_addr_U <= pix_y(5 downto 0) - U_y_t_u(5 downto 0);
    rom_col_U <= pix_x(5 downto 0) - U_x_l_u(5 downto 0);
    rom_data_U <= U_ROM(to_integer(rom_addr_U));
    rom_bit_U <= rom_data_U(to_integer(rom_col_U));

    
    rom_addr_D_1 <= pix_y(5 downto 0) - D_1_y_t_u(5 downto 0);
    rom_col_D_1 <= pix_x(5 downto 0) - D_1_x_l_u(5 downto 0);
    rom_data_D_1 <= D_1_ROM(to_integer(rom_addr_D_1));
    rom_bit_D_1 <= rom_data_D_1(to_integer(rom_col_D_1));

    
    rom_addr_I <= pix_y(5 downto 0) - I_y_t_u(5 downto 0);
    rom_col_I <= pix_x(5 downto 0) - I_x_l_u(5 downto 0);
    rom_data_I <= I_ROM(to_integer(rom_addr_I));
    rom_bit_I <= rom_data_I(to_integer(rom_col_I));

    
    rom_addr_E <= pix_y(5 downto 0) - E_y_t_u(5 downto 0);
    rom_col_E <= pix_x(5 downto 0) - E_x_l_u(5 downto 0);
    rom_data_E <= E_ROM(to_integer(rom_addr_E));
    rom_bit_E <= rom_data_E(to_integer(rom_col_E));

    
    rom_addr_D_2 <= pix_y(5 downto 0) - D_2_y_t_u(5 downto 0);
    rom_col_D_2 <= pix_x(5 downto 0) - D_2_x_l_u(5 downto 0);
    rom_data_D_2 <= D_2_ROM(to_integer(rom_addr_D_2));
    rom_bit_D_2 <= rom_data_D_2(to_integer(rom_col_D_2));

    U_cur_val_on <= '1' when (sq_U_on = '1') and (rom_bit_U = '1') and (life_cnter = "00") else '0';
    D_1_cur_val_on <= '1' when (sq_D_1_on = '1') and (rom_bit_D_1 = '1') and (life_cnter = "00") else '0';
    I_cur_val_on <= '1' when (sq_I_on = '1') and (rom_bit_I = '1') and (life_cnter = "00") else '0';
    E_cur_val_on <= '1' when (sq_E_on = '1') and (rom_bit_E = '1') and (life_cnter = "00") else '0';
    D_2_cur_val_on <= '1' when (sq_D_2_on = '1') and (rom_bit_D_2 = '1') and (life_cnter = "00") else '0';

    graph_rgb <= char_rgb when U_cur_val_on = '1' else 
        char_rgb when D_1_cur_val_on = '1' else
        char_rgb when I_cur_val_on = '1' else
        char_rgb when E_cur_val_on = '1' else
        char_rgb when D_2_cur_val_on = '1' else
        "000";
    
    game_over_on <= '1' when (life_cnter = "00") else '0';
end arch;